
module  ALU(
    input A,
    input B,
    input operator,
    output carry,
    output overflow,
    output result,
    output zero
);
//add:000

//sub:001

//shift

//compare

//judge:overflow/C/O


endmodule // ALU
